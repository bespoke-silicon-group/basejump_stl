module basic_checker
  import bsg_cache_pkg::*;
  #(parameter data_width_p="inv"
    , parameter addr_width_p="inv"
    , parameter mem_size_p="inv"

    , parameter data_mask_width_lp=(data_width_p>>3)
    , parameter cache_pkt_width_lp= `bsg_cache_pkt_width(addr_width_p,data_width_p)
  ) 
  (
    input clk_i
    , input reset_i
      
    , input en_i

    , input [cache_pkt_width_lp-1:0] cache_pkt_i
    , input v_i
    , input ready_o

    , input [data_width_p-1:0] data_o
    , input v_o
    , input yumi_i
  );


  `declare_bsg_cache_pkt_s(addr_width_p,data_width_p);

  bsg_cache_pkt_s cache_pkt;
  assign cache_pkt = cache_pkt_i;

  logic [data_width_p-1:0] shadow_mem [mem_size_p-1:0];
  logic [data_width_p-1:0] result [*];

  wire [addr_width_p-1:0] cache_pkt_word_addr = cache_pkt.addr[addr_width_p-1:3];

  // store logic
  logic [data_width_p-1:0] load_data, load_data_final;
  logic [data_width_p-1:0] store_pre_data;
  logic [data_width_p-1:0] store_data;
  logic [data_mask_width_lp-1:0] store_mask;

  always_comb begin
    case (cache_pkt.opcode)
      AMOOR_D, AMOOR_W: begin
        store_pre_data = cache_pkt.data | load_data_final;
      end
      default: begin
        store_pre_data = cache_pkt.data;
      end
    endcase
  end

  always_comb begin
    case (cache_pkt.opcode)
      
      SD, AMOSWAP_D, AMOOR_D: begin
        store_data = store_pre_data;
        store_mask = 8'b1111_1111;
      end

      SW, AMOSWAP_W, AMOOR_W: begin
        store_data = {2{store_pre_data[31:0]}};
        store_mask = {
          {4{ cache_pkt.addr[2]}},
          {4{~cache_pkt.addr[2]}}
        };
      end

      SH: begin
        store_data = {4{store_pre_data[15:0]}};
        store_mask = {
          {2{ cache_pkt.addr[2] &  cache_pkt.addr[1]}},
          {2{ cache_pkt.addr[2] & ~cache_pkt.addr[1]}},
          {2{~cache_pkt.addr[2] &  cache_pkt.addr[1]}},
          {2{~cache_pkt.addr[2] & ~cache_pkt.addr[1]}}
        };
      end

      SB: begin
        store_data = {8{store_pre_data[7:0]}};
        store_mask = {
           { cache_pkt.addr[2] &  cache_pkt.addr[1] &   cache_pkt.addr[0]},
           { cache_pkt.addr[2] &  cache_pkt.addr[1] &  ~cache_pkt.addr[0]},
           { cache_pkt.addr[2] & ~cache_pkt.addr[1] &   cache_pkt.addr[0]},
           { cache_pkt.addr[2] & ~cache_pkt.addr[1] &  ~cache_pkt.addr[0]},
           {~cache_pkt.addr[2] &  cache_pkt.addr[1] &   cache_pkt.addr[0]},
           {~cache_pkt.addr[2] &  cache_pkt.addr[1] &  ~cache_pkt.addr[0]},
           {~cache_pkt.addr[2] & ~cache_pkt.addr[1] &   cache_pkt.addr[0]},
           {~cache_pkt.addr[2] & ~cache_pkt.addr[1] &  ~cache_pkt.addr[0]}
        };
      end

      SM: begin
        store_data = store_pre_data;
        store_mask = cache_pkt.mask;
      end

      default: begin
        store_data = '0;
        store_mask = '0;
      end
    endcase
  end

  // load logic
  logic [7:0] byte_sel;
  logic [15:0] half_sel;
  logic [31:0] word_sel;

  assign load_data = shadow_mem[cache_pkt_word_addr];

  bsg_mux #(
    .els_p(8)
    ,.width_p(8)
  ) byte_mux (
    .data_i(load_data)
    ,.sel_i(cache_pkt.addr[2:0])
    ,.data_o(byte_sel)
  );

  bsg_mux #(
    .els_p(4)
    ,.width_p(16)
  ) half_mux (
    .data_i(load_data)
    ,.sel_i(cache_pkt.addr[2:1])
    ,.data_o(half_sel)
  );

  bsg_mux #(
    .els_p(2)
    ,.width_p(32)
  ) word_mux (
    .data_i(load_data)
    ,.sel_i(cache_pkt.addr[2])
    ,.data_o(word_sel)
  );


  always_comb begin
    case (cache_pkt.opcode)
      LD, AMOSWAP_D, AMOOR_D: load_data_final = load_data;
      LW, AMOSWAP_W, AMOOR_W: load_data_final = {{32{word_sel[31]}}, word_sel};
      LH: load_data_final = {{48{half_sel[15]}}, half_sel};
      LB: load_data_final = {{56{byte_sel[7]}}, byte_sel};
      LWU: load_data_final = {{32{1'b0}}, word_sel};
      LHU: load_data_final = {{48{1'b0}}, half_sel};
      LBU: load_data_final = {{56{1'b0}}, byte_sel};
      default: load_data_final = '0;
    endcase
  end



  integer send_id, recv_id;

  always_ff @ (posedge clk_i) begin
    if (reset_i) begin
      send_id <= '0;
      recv_id <= '0;
      for (integer i = 0; i < mem_size_p; i++)
        shadow_mem[i] = '0;
    end
    else begin

      if (en_i) begin

        // input recorder
        if (v_i & ready_o) begin
          case (cache_pkt.opcode)

            TAGST: begin
              result[send_id] = '0;
              send_id++;
            end

            LD, LW, LH, LB, LWU, LHU, LBU: begin
              result[send_id] = load_data_final;
              send_id++;
            end

            SD, SW, SH, SB: begin
              result[send_id] = '0;
              send_id++;
              for (integer i = 0; i < data_mask_width_lp; i++)
                if (store_mask[i])
                  shadow_mem[cache_pkt_word_addr][8*i+:8] <= store_data[8*i+:8];
            end

            AMOSWAP_W, AMOOR_W,
            AMOSWAP_D, AMOOR_D: begin
              result[send_id] = load_data_final;
              send_id++;
              for (integer i = 0; i < data_mask_width_lp; i++)
                if (store_mask[i])
                  shadow_mem[cache_pkt_word_addr][8*i+:8] <= store_data[8*i+:8];
            end

          endcase
        end

        // output checker
        if (v_o & yumi_i) begin
          assert(result[recv_id] == data_o)
            else $fatal("[BSG_FATAL] output does not match expected result. Id=%d, Expected: %x. Actual: %x.",
                    recv_id, result[recv_id], data_o);
          recv_id++;
        end
      end
    end
  end

  
endmodule
