//File contains list of macros used in the DMC testbench.

`define bsg_log_utils(ARG) \
	string msg_id = ``ARG;
