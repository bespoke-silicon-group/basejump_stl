`include "bsg_defines.sv"

module bsg_clkinv #(parameter width_p=1
                    , parameter strength_p=8
                    , parameter harden_p=0
                    )
   (input    [width_p-1:0] i
    , output [width_p-1:0] o
    );

   assign o = ~i;

endmodule
