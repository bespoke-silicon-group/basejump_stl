//TODO: akashs3: why are these defines? why not enums?
`define WRITE 3'b000
`define READ  3'b001
