package bsg_dmc_tests_pkg;
	import uvm_pkg::*;
	import bsg_dmc_pkg::*;
	import bsg_dmc_asic_pkg::*;

	`include "../env/bsg_dmc_env.sv"
	`include "bsg_dmc_base_test.sv"
endpackage
