interface bsg_dmc_ddr_interface;

