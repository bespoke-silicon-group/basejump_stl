interface bsg_dmc_dfi_interface;
	logic                          	dfi_clk_1x_i;
	logic                          	dfi_clk_2x_i;
	logic                          	dfi_rst_i;
	logic                    [2:0] 	dfi_bank_i;
	logic                   [15:0] 	dfi_address_i;
	logic                          	dfi_cke_i;
	logic                          	dfi_cs_n_i;
	logic                          	dfi_ras_n_i;
	logic                          	dfi_cas_n_i;
	logic                          	dfi_we_n_i;
	logic                          	dfi_reset_n_i;
	logic                          	dfi_odt_i;
	logic                          	dfi_wrdata_en_i;
	logic  [2*dq_data_width_p-1:0] 	dfi_wrdata_i;
	logic      [2*dq_group_lp-1:0] 	dfi_wrdata_mask_i;
	logic                          	dfi_rddata_en_i;
	logic [2*dq_data_width_p-1:0] 	dfi_rddata_o;
	logic                   		dfi_rddata_valid_o;
endinterface
