package bsg_dmc_seq_pkg;
	import uvm_pkg::*;
	import bsg_dmc_pkg::*;
	import bsg_dmc_asic_pkg::*;
	import bsg_dmc_params_pkg::*;
	
	`include "bsg_dmc_cmd_seq.sv"
	`include "bsg_dmc_write_seq.sv"
	`include "bsg_dmc_read_seq.sv"
	`include "bsg_dmc_top_seq.sv"

endpackage: bsg_dmc_seq_pkg
