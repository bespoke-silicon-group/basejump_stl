module test_bsg
#(parameter num_out_p=-1,
  parameter cycle_time_p=10,
  parameter reset_cycles_lo_p=-1,
  parameter reset_cycles_hi_p=-1
  );

  wire clk;
  wire reset;

  bsg_nonsynth_clock_gen #(  .cycle_time_p(cycle_time_p)
                          )  clock_gen
                          (  .o(clk)
                          );

  bsg_nonsynth_reset_gen #(  .num_clocks_p     (1)
                           , .reset_cycles_lo_p(reset_cycles_lo_p)
                           , .reset_cycles_hi_p(reset_cycles_hi_p)
                          )  reset_gen
                          (  .clk_i        (clk) 
                           , .async_reset_o(reset)
                          );

  initial begin
    $display("[BSG_PASS] Empty testbench");
    $finish();
  end
  
  wire [`BSG_SAFE_CLOG2(num_out_p)-1:0] i;
  wire v_i;
  wire [num_out_p-1:0] o;

  bsg_decode_with_v #(
    .num_out_p(num_out_p))
    DUT (
    .i(i),
    .v_i(v_i),
    .o(o)
  );

endmodule
