/**
 *  bsg_cache_non_blocking_tl_stage.v
 *
 *  tag-lookup stage
 *
 *  @author tommy
 *
 */



module bsg_cache_non_blocking_tl_stage
  #(
  )
  (
    input clk_i
    , input reset_i

    
  );




endmodule
