package bsg_dmc_params_pkg;

	`include "bsg_dmc_defines.vh"
	`include "bsg_dmc_params.vh"

endpackage: bsg_dmc_params_pkg
