/**
 *    bsg_cache_non_blocking_stat_mem.v
 *
 *    stat_mem and peripheral circuits
 *
 *    @author tommy
 *
 */


module bsg_cache_non_blocking_stat_mem
  #(parameter ways_p="inv"
    , parameter sets_p="inv"
  )
  (
    input clk_i
    , input reset_i

  );





endmodule
