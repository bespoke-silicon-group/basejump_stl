package bsg_dmc_params_pkg;

	`include "bsg_dmc_defines.vh"
	`include "bsg_dmc_params.vh"
	`include "bsg_dmc_macros.sv"

endpackage: bsg_dmc_params_pkg
