module bsg_nonsynth_random_yumi_gen 
  #(parameter `BSG_INV_PARAM(yumi_min_delay_p)
    , parameter `BSG_INV_PARAM(yumi_max_delay_p)
  )
  (
    input clk_i
    , input reset_i
    
    , input v_i
    , output logic yumi_o
  );


  integer yumi_count_r;
  
  always_ff @ (posedge clk_i) begin
    if (reset_i) begin
      yumi_count_r <= $urandom() % (yumi_max_delay_p-yumi_min_delay_p) + yumi_min_delay_p;
    end
    else begin
      if (v_i) begin
        if (yumi_count_r <= 0) begin
          yumi_count_r <= $urandom() % (yumi_max_delay_p-yumi_min_delay_p) + yumi_min_delay_p;
        end
        else begin
          yumi_count_r <= yumi_count_r - 1;
        end
      end
    end
  end

  assign yumi_o = v_i & (yumi_count_r == 0);
  

endmodule

`BSG_ABSTRACT_MODULE(bsg_nonsynth_random_yumi_gen)
