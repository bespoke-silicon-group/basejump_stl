
  module bsg_mem_1r1w_sync_w64_d512_m2_hard;
      bsg_mem_1r1w_sync_synth #(
        .width_p(64)
        ,.els_p(512)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1r1w_sync_w32_d1024_m2_hard;
      bsg_mem_1r1w_sync_synth #(
        .width_p(32)
        ,.els_p(1024)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1r1w_sync_mask_write_bit_w64_d512_m2_hard;
      bsg_mem_1r1w_sync_mask_write_bit_synth #(
        .width_p(64)
        ,.els_p(512)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1r1w_sync_mask_write_bit_w32_d1024_m2_hard;
      bsg_mem_1r1w_sync_mask_write_bit_synth #(
        .width_p(32)
        ,.els_p(1024)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1r1w_sync_mask_write_byte_w64_d512_m2_hard;
      bsg_mem_1r1w_sync_mask_write_byte_synth #(
        .width_p(64)
        ,.els_p(512)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1r1w_sync_mask_write_byte_w32_d1024_m2_hard;
      bsg_mem_1r1w_sync_mask_write_byte_synth #(
        .width_p(32)
        ,.els_p(1024)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1rw_sync_w64_d512_m2_hard;
      bsg_mem_1rw_sync_synth #(
        .width_p(64)
        ,.els_p(512)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1rw_sync_w32_d128_m2_hard;
      bsg_mem_1rw_sync_synth #(
        .width_p(32)
        ,.els_p(128)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1rw_sync_mask_write_bit_w64_d512_m2_hard;
      bsg_mem_1rw_sync_mask_write_bit_synth #(
        .width_p(64)
        ,.els_p(512)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1rw_sync_mask_write_bit_w32_d128_m2_hard;
      bsg_mem_1rw_sync_mask_write_bit_synth #(
        .width_p(32)
        ,.els_p(128)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1rw_sync_mask_write_byte_w64_d512_m2_hard;
      bsg_mem_1rw_sync_mask_write_byte_synth #(
        .width_p(64)
        ,.els_p(512)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_1rw_sync_mask_write_byte_w32_d128_m2_hard;
      bsg_mem_1rw_sync_mask_write_byte_synth #(
        .width_p(32)
        ,.els_p(128)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_2r1w_sync_w64_d32_m2_hard;
      bsg_mem_2r1w_sync_synth #(
        .width_p(64)
        ,.els_p(32)
      ) func (.*);
  endmodule
  
  

  module bsg_mem_3r1w_sync_w66_d32_m2_hard;
      bsg_mem_3r1w_sync_synth #(
        .width_p(66)
        ,.els_p(32)
      ) func (.*);
  endmodule
  
  
