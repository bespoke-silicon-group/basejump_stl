///////////////////////////////////////////////////////////////////////////////////////////////////
//    		BASEJUMP STL
//
//       MODULE: bsg_dmc_trace_to_xilinx_ui_adapter
//  DESCRIPTION: Takes the DMC cmd, addr, wdata, wmask trace packet and converts into XILINX UI interface to feed to DMC;
//  			 And converts UI read interface signals to trace packet to forward to FPGA
//    AUTHOR(S): Akash Suresh, akashs3@uw.edu
// ORGANIZATION: Bespoke Silicon Group, University of Washington
//      CREATED: 01/07/22
///////////////////////////////////////////////////////////////////////////////////////////////////
module bsg_dmc_trace_to_xilinx_ui_adapter
	import bsg_dmc_pkg::*;
	#(	parameter `BSG_INV_PARAM( data_width_p),
		parameter `BSG_INV_PARAM( addr_width_p),
		parameter `BSG_INV_PARAM( cmd_width_p),
		parameter `BSG_INV_PARAM( burst_width_p),

		localparam payload_width_lp = data_width_p + (data_width_p>>3) + 4,
		localparam mask_width_lp = data_width_p>>3,
        localparam read_data_buffer_size_lp = burst_width_p*2
	)
	( 	input 									core_clk_i,
		input									core_reset_i,

        // Trace data from producer
		output      							ready_o,
		input [payload_width_lp -1 :0] 			data_i,
		input 									v_i,

        // Read data to consumer
		output logic [data_width_p -1 :0]	    data_o,
		output logic							v_o,
        input                                   yumi_i,

   		// xilinx user interface
   		output logic [addr_width_p-1:0]        	app_addr_o,
   		output app_cmd_e				    	app_cmd_o,
   		output logic                       		app_en_o,
   		input                              		app_rdy_i,
   		output logic                       		app_wdf_wren_o,
   		output logic [data_width_p-1:0]			app_wdf_data_o,
   		output logic [(data_width_p>>3)-1:0] 	app_wdf_mask_o,
   		output logic                   			app_wdf_end_o,
   		input                              		app_wdf_rdy_i,
   		input                              		app_rd_data_valid_i,
   		input [data_width_p-1:0] 		      	app_rd_data_i,
   		input                              		app_rd_data_end_i
	);

    localparam cmd_trace_zero_padding_width_lp = data_width_p + mask_width_lp - cmd_width_p - addr_width_p;
	`declare_dmc_cmd_trace_entry_s(addr_width_p, cmd_trace_zero_padding_width_lp)
	`declare_dmc_wdata_trace_entry_s(data_width_p, mask_width_lp)

	// counter to load one packet per burst per cycle onto app_wdata and app_wmask
	logic [`BSG_SAFE_CLOG2(burst_width_p) - 1:0] write_count;

	logic burst_done;
    logic read_data_valid_li, read_data_fifo_ready_lo;
    logic [`BSG_SAFE_CLOG2(read_data_buffer_size_lp) -1 :0] read_credit;

	dmc_cmd_trace_entry_s cmd_trace_data;
	dmc_data_trace_entry_s wdata_trace_data;

	assign cmd_trace_data = data_i;
    assign wdata_trace_data = data_i;

	assign ready_o =  app_rdy_i;

	assign burst_done =  (write_count == burst_width_p  - 1);

	assign is_write = (v_i && cmd_trace_data.cmd_wdata_n) ? ((cmd_trace_data.cmd == WP) || (cmd_trace_data.cmd == WR) )  : 0;

	assign app_wdf_end_o = burst_done & app_wdf_wren_o;

	assign {feed_to_app_wdata, feed_to_app_wmask} = data_i;
	
	// counting write_count per burst
	bsg_counter_clear_up
					#(.max_val_p(burst_width_p - 1)
					,.init_val_p(0)
                    ,.disable_overflow_warning_p(1))
					write_counter
					(.clk_i(core_clk_i)
					,.reset_i(core_reset_i)
					,.clear_i(1'b0)                        
					,.up_i(app_wdf_wren_o & app_wdf_rdy_i )
					,.count_o(write_count)
					);
	
	// Convert UI command and addr
    always_comb begin
        if(v_i &&   app_rdy_i && cmd_trace_data.cmd_wdata_n ) begin
            if((cmd_trace_data.cmd == WR) || (cmd_trace_data.cmd == WP) && app_wdf_rdy_i) begin
                app_en_o = 1;
            end
            else if((cmd_trace_data.cmd == RD) || (cmd_trace_data.cmd == RP) && (read_credit >= burst_width_p)) begin
                app_en_o = 1;
            end
        end
        else begin
            app_en_o = 0;
        end
    end

	assign app_cmd_o = cmd_trace_data.cmd;
	assign app_addr_o = cmd_trace_data.addr;

    always @(posedge core_clk_i) begin
        if(core_reset_i) begin
            app_wdf_wren_o <= 0;
        end
        else if(is_write && app_wdf_rdy_i & v_i) begin
            app_wdf_wren_o <= 1;
        end
        else if(burst_done) begin
            app_wdf_wren_o <= 0;
        end
    end

    assign app_wdf_data_o = wdata_trace_data.data;
    assign app_wdf_mask_o = wdata_trace_data.mask;

    assign read_data_valid_li = app_rd_data_valid_i & read_data_fifo_ready_lo; 

    bsg_fifo_1r1w_small 
    				#(.width_p(data_width_p)
    				,.els_p(read_data_buffer_size_lp)
    				) read_data_fifo
    				(.clk_i  (core_clk_i)
    				,.reset_i(core_reset_i)
    				
    				,.ready_o(read_data_fifo_ready_lo)
    				,.data_i (app_rd_data_i)
    				,.v_i    (app_rd_data_valid_i)
    				
    				,.v_o    (v_o)
    				,.data_o (data_o)
    				,.yumi_i (v_o & yumi_i)
    				);

    always@(posedge core_clk_i) begin
        if(core_reset_i) begin
            read_credit <= read_data_buffer_size_lp -1 ;
        end
        if(app_rd_data_valid_i && !app_rd_data_end_i) begin
            read_credit <= read_credit - 1;
        end
        else if(app_rd_data_end_i) begin
            read_credit <= read_credit + burst_width_p - 1;
        end
    end

endmodule
