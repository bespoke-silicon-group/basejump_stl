module bsg_mesosync_io()











endmodule
